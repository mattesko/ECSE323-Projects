library verilog;
use verilog.vl_types.all;
entity testing2_vlg_vec_tst is
end testing2_vlg_vec_tst;
