library verilog;
use verilog.vl_types.all;
entity g27_dealer_vlg_vec_tst is
end g27_dealer_vlg_vec_tst;
