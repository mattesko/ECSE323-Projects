library verilog;
use verilog.vl_types.all;
entity g27_modulo_vlg_vec_tst is
end g27_modulo_vlg_vec_tst;
