library verilog;
use verilog.vl_types.all;
entity g27_shift_left_3_vlg_vec_tst is
end g27_shift_left_3_vlg_vec_tst;
