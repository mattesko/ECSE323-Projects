library ieee;
use ieee.std_logic_1164.all;

entity p_enable is
	port(addr : in std_logic_vector(5 downto 0);
		  p_en : out std_logic_vector(51 downto 0));
end p_enable;

architecture p_enable_arch of p_enable is
begin
with addr select p_en <=
"1111111111111111111111111111111111111111111111111111" when "000000",
"1111111111111111111111111111111111111111111111111110" when "000001",
"1111111111111111111111111111111111111111111111111100" when "000010",
"1111111111111111111111111111111111111111111111111000" when "000011",
"1111111111111111111111111111111111111111111111110000" when "000100",
"1111111111111111111111111111111111111111111111100000" when "000101",
"1111111111111111111111111111111111111111111111000000" when "000110",
"1111111111111111111111111111111111111111111110000000" when "000111",
"1111111111111111111111111111111111111111111100000000" when "001000",
"1111111111111111111111111111111111111111111000000000" when "001001",
"1111111111111111111111111111111111111111110000000000" when "001010",
"1111111111111111111111111111111111111111100000000000" when "001011",
"1111111111111111111111111111111111111111000000000000" when "001100",
"1111111111111111111111111111111111111110000000000000" when "001101",
"1111111111111111111111111111111111111100000000000000" when "001110",
"1111111111111111111111111111111111111000000000000000" when "001111",
"1111111111111111111111111111111111110000000000000000" when "010000",
"1111111111111111111111111111111111100000000000000000" when "010001",
"1111111111111111111111111111111111000000000000000000" when "010010",
"1111111111111111111111111111111110000000000000000000" when "010011",
"1111111111111111111111111111111100000000000000000000" when "010100",
"1111111111111111111111111111111000000000000000000000" when "010101",
"1111111111111111111111111111110000000000000000000000" when "010110",
"1111111111111111111111111111100000000000000000000000" when "010111",
"1111111111111111111111111111000000000000000000000000" when "011000",
"1111111111111111111111111110000000000000000000000000" when "011001",
"1111111111111111111111111100000000000000000000000000" when "011010",
"1111111111111111111111111000000000000000000000000000" when "011011",
"1111111111111111111111110000000000000000000000000000" when "011100",
"1111111111111111111111100000000000000000000000000000" when "011101",
"1111111111111111111111000000000000000000000000000000" when "011110",
"1111111111111111111110000000000000000000000000000000" when "011111",
"1111111111111111111100000000000000000000000000000000" when "100000",
"1111111111111111111000000000000000000000000000000000" when "100001",
"1111111111111111110000000000000000000000000000000000" when "100010",
"1111111111111111100000000000000000000000000000000000" when "100011",
"1111111111111111000000000000000000000000000000000000" when "100100",
"1111111111111110000000000000000000000000000000000000" when "100101",
"1111111111111100000000000000000000000000000000000000" when "100110",
"1111111111111000000000000000000000000000000000000000" when "100111",
"1111111111110000000000000000000000000000000000000000" when "101000",
"1111111111100000000000000000000000000000000000000000" when "101001",
"1111111111000000000000000000000000000000000000000000" when "101010",
"1111111110000000000000000000000000000000000000000000" when "101011",
"1111111100000000000000000000000000000000000000000000" when "101100",
"1111111000000000000000000000000000000000000000000000" when "101101",
"1111110000000000000000000000000000000000000000000000" when "101110",
"1111100000000000000000000000000000000000000000000000" when "101111",
"1111000000000000000000000000000000000000000000000000" when "110000",
"1110000000000000000000000000000000000000000000000000" when "110001",
"1100000000000000000000000000000000000000000000000000" when "110010",
"1000000000000000000000000000000000000000000000000000" when "110011",
"0000000000000000000000000000000000000000000000000000" when others;
end;
	