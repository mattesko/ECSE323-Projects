library verilog;
use verilog.vl_types.all;
entity g27_decision_maker_FSM_schematic_vlg_vec_tst is
end g27_decision_maker_FSM_schematic_vlg_vec_tst;
