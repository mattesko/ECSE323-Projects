library verilog;
use verilog.vl_types.all;
entity g27_lab1_vlg_check_tst is
    port(
        AeqB            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g27_lab1_vlg_check_tst;
