library verilog;
use verilog.vl_types.all;
entity rand_modulo_test_vlg_vec_tst is
end rand_modulo_test_vlg_vec_tst;
