library verilog;
use verilog.vl_types.all;
entity g27_6bit_shift_right_matthew_vlg_vec_tst is
end g27_6bit_shift_right_matthew_vlg_vec_tst;
