library verilog;
use verilog.vl_types.all;
entity g27_lab1_vlg_vec_tst is
end g27_lab1_vlg_vec_tst;
