-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Nov 01 22:31:02 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY g27_stack52 IS 
	PORT
	(
		ENABLE :  IN  STD_LOGIC;
		RST :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		ADDR :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		DATA :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		MODE :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		EMPTY :  OUT  STD_LOGIC;
		PUSH :  OUT  STD_LOGIC;
		POP :  OUT  STD_LOGIC;
		FULL :  OUT  STD_LOGIC;
		NUM :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		VALUE :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END g27_stack52;

ARCHITECTURE bdf_type OF g27_stack52 IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT lpm_ff_0
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_0: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_0: COMPONENT IS true;

COMPONENT lpm_ff_1
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_1: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_1: COMPONENT IS true;

COMPONENT lpm_ff_12
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_12: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_12: COMPONENT IS true;

COMPONENT lpm_ff_14
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_14: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_14: COMPONENT IS true;

COMPONENT lpm_ff_16
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_16: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_16: COMPONENT IS true;

COMPONENT lpm_ff_18
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_18: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_18: COMPONENT IS true;

COMPONENT lpm_ff_2
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_2: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_2: COMPONENT IS true;

COMPONENT lpm_ff_20
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_20: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_20: COMPONENT IS true;

COMPONENT lpm_ff_3
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_3: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_3: COMPONENT IS true;

COMPONENT lpm_ff_5
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_5: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_5: COMPONENT IS true;

COMPONENT lpm_ff_7
	PORT(enable : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 sclr : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ff_7: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ff_7: COMPONENT IS true;

TYPE ARRAY2D0 IS ARRAY (51 DOWNTO 0,5 DOWNTO 0) OF STD_LOGIC;

COMPONENT lpm_mux_6
	PORT(data : IN ARRAY2D0;
		 sel : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
END COMPONENT;
ATTRIBUTE black_box OF lpm_mux_6: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_mux_6: COMPONENT IS true;

COMPONENT busmux_10
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_10: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_10: COMPONENT IS true;

COMPONENT busmux_11
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_11: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_11: COMPONENT IS true;

COMPONENT busmux_13
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_13: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_13: COMPONENT IS true;

COMPONENT busmux_15
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_15: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_15: COMPONENT IS true;

COMPONENT busmux_17
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_17: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_17: COMPONENT IS true;

COMPONENT busmux_19
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_19: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_19: COMPONENT IS true;

COMPONENT busmux_21
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_21: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_21: COMPONENT IS true;

COMPONENT busmux_22
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_22: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_22: COMPONENT IS true;

COMPONENT busmux_4
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_4: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_4: COMPONENT IS true;

COMPONENT busmux_8
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_8: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_8: COMPONENT IS true;

COMPONENT busmux_9
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_9: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_9: COMPONENT IS true;

COMPONENT lpm_counter0
	PORT(sclr : IN STD_LOGIC;
		 sload : IN STD_LOGIC;
		 sset : IN STD_LOGIC;
		 updown : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 cnt_en : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux2
	PORT(data0x : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT g27_pop_enable
	PORT(clk : IN STD_LOGIC;
		 N : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 P_EN : OUT STD_LOGIC_VECTOR(51 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	0 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	10 :  STD_LOGIC;
SIGNAL	100 :  STD_LOGIC;
SIGNAL	101 :  STD_LOGIC;
SIGNAL	102 :  STD_LOGIC;
SIGNAL	103 :  STD_LOGIC;
SIGNAL	104 :  STD_LOGIC;
SIGNAL	105 :  STD_LOGIC;
SIGNAL	11 :  STD_LOGIC;
SIGNAL	110 :  STD_LOGIC;
SIGNAL	111 :  STD_LOGIC;
SIGNAL	112 :  STD_LOGIC;
SIGNAL	113 :  STD_LOGIC;
SIGNAL	114 :  STD_LOGIC;
SIGNAL	115 :  STD_LOGIC;
SIGNAL	12 :  STD_LOGIC;
SIGNAL	120 :  STD_LOGIC;
SIGNAL	121 :  STD_LOGIC;
SIGNAL	122 :  STD_LOGIC;
SIGNAL	123 :  STD_LOGIC;
SIGNAL	124 :  STD_LOGIC;
SIGNAL	125 :  STD_LOGIC;
SIGNAL	13 :  STD_LOGIC;
SIGNAL	130 :  STD_LOGIC;
SIGNAL	131 :  STD_LOGIC;
SIGNAL	132 :  STD_LOGIC;
SIGNAL	133 :  STD_LOGIC;
SIGNAL	134 :  STD_LOGIC;
SIGNAL	135 :  STD_LOGIC;
SIGNAL	14 :  STD_LOGIC;
SIGNAL	140 :  STD_LOGIC;
SIGNAL	141 :  STD_LOGIC;
SIGNAL	142 :  STD_LOGIC;
SIGNAL	143 :  STD_LOGIC;
SIGNAL	144 :  STD_LOGIC;
SIGNAL	145 :  STD_LOGIC;
SIGNAL	15 :  STD_LOGIC;
SIGNAL	150 :  STD_LOGIC;
SIGNAL	151 :  STD_LOGIC;
SIGNAL	152 :  STD_LOGIC;
SIGNAL	153 :  STD_LOGIC;
SIGNAL	154 :  STD_LOGIC;
SIGNAL	155 :  STD_LOGIC;
SIGNAL	16 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	17 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	18 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	19 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	20 :  STD_LOGIC;
SIGNAL	200 :  STD_LOGIC;
SIGNAL	201 :  STD_LOGIC;
SIGNAL	202 :  STD_LOGIC;
SIGNAL	203 :  STD_LOGIC;
SIGNAL	204 :  STD_LOGIC;
SIGNAL	205 :  STD_LOGIC;
SIGNAL	21 :  STD_LOGIC;
SIGNAL	210 :  STD_LOGIC;
SIGNAL	211 :  STD_LOGIC;
SIGNAL	212 :  STD_LOGIC;
SIGNAL	213 :  STD_LOGIC;
SIGNAL	214 :  STD_LOGIC;
SIGNAL	215 :  STD_LOGIC;
SIGNAL	22 :  STD_LOGIC;
SIGNAL	220 :  STD_LOGIC;
SIGNAL	221 :  STD_LOGIC;
SIGNAL	222 :  STD_LOGIC;
SIGNAL	223 :  STD_LOGIC;
SIGNAL	224 :  STD_LOGIC;
SIGNAL	225 :  STD_LOGIC;
SIGNAL	23 :  STD_LOGIC;
SIGNAL	230 :  STD_LOGIC;
SIGNAL	231 :  STD_LOGIC;
SIGNAL	232 :  STD_LOGIC;
SIGNAL	233 :  STD_LOGIC;
SIGNAL	234 :  STD_LOGIC;
SIGNAL	235 :  STD_LOGIC;
SIGNAL	24 :  STD_LOGIC;
SIGNAL	240 :  STD_LOGIC;
SIGNAL	241 :  STD_LOGIC;
SIGNAL	242 :  STD_LOGIC;
SIGNAL	243 :  STD_LOGIC;
SIGNAL	244 :  STD_LOGIC;
SIGNAL	245 :  STD_LOGIC;
SIGNAL	25 :  STD_LOGIC;
SIGNAL	250 :  STD_LOGIC;
SIGNAL	251 :  STD_LOGIC;
SIGNAL	252 :  STD_LOGIC;
SIGNAL	253 :  STD_LOGIC;
SIGNAL	254 :  STD_LOGIC;
SIGNAL	255 :  STD_LOGIC;
SIGNAL	26 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	27 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	28 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	29 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	30 :  STD_LOGIC;
SIGNAL	300 :  STD_LOGIC;
SIGNAL	301 :  STD_LOGIC;
SIGNAL	302 :  STD_LOGIC;
SIGNAL	303 :  STD_LOGIC;
SIGNAL	304 :  STD_LOGIC;
SIGNAL	305 :  STD_LOGIC;
SIGNAL	31 :  STD_LOGIC;
SIGNAL	310 :  STD_LOGIC;
SIGNAL	311 :  STD_LOGIC;
SIGNAL	312 :  STD_LOGIC;
SIGNAL	313 :  STD_LOGIC;
SIGNAL	314 :  STD_LOGIC;
SIGNAL	315 :  STD_LOGIC;
SIGNAL	32 :  STD_LOGIC;
SIGNAL	320 :  STD_LOGIC;
SIGNAL	321 :  STD_LOGIC;
SIGNAL	322 :  STD_LOGIC;
SIGNAL	323 :  STD_LOGIC;
SIGNAL	324 :  STD_LOGIC;
SIGNAL	325 :  STD_LOGIC;
SIGNAL	33 :  STD_LOGIC;
SIGNAL	330 :  STD_LOGIC;
SIGNAL	331 :  STD_LOGIC;
SIGNAL	332 :  STD_LOGIC;
SIGNAL	333 :  STD_LOGIC;
SIGNAL	334 :  STD_LOGIC;
SIGNAL	335 :  STD_LOGIC;
SIGNAL	34 :  STD_LOGIC;
SIGNAL	340 :  STD_LOGIC;
SIGNAL	341 :  STD_LOGIC;
SIGNAL	342 :  STD_LOGIC;
SIGNAL	343 :  STD_LOGIC;
SIGNAL	344 :  STD_LOGIC;
SIGNAL	345 :  STD_LOGIC;
SIGNAL	35 :  STD_LOGIC;
SIGNAL	350 :  STD_LOGIC;
SIGNAL	351 :  STD_LOGIC;
SIGNAL	352 :  STD_LOGIC;
SIGNAL	353 :  STD_LOGIC;
SIGNAL	354 :  STD_LOGIC;
SIGNAL	355 :  STD_LOGIC;
SIGNAL	36 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	37 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	38 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	39 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	40 :  STD_LOGIC;
SIGNAL	400 :  STD_LOGIC;
SIGNAL	401 :  STD_LOGIC;
SIGNAL	402 :  STD_LOGIC;
SIGNAL	403 :  STD_LOGIC;
SIGNAL	404 :  STD_LOGIC;
SIGNAL	405 :  STD_LOGIC;
SIGNAL	41 :  STD_LOGIC;
SIGNAL	410 :  STD_LOGIC;
SIGNAL	411 :  STD_LOGIC;
SIGNAL	412 :  STD_LOGIC;
SIGNAL	413 :  STD_LOGIC;
SIGNAL	414 :  STD_LOGIC;
SIGNAL	415 :  STD_LOGIC;
SIGNAL	42 :  STD_LOGIC;
SIGNAL	420 :  STD_LOGIC;
SIGNAL	421 :  STD_LOGIC;
SIGNAL	422 :  STD_LOGIC;
SIGNAL	423 :  STD_LOGIC;
SIGNAL	424 :  STD_LOGIC;
SIGNAL	425 :  STD_LOGIC;
SIGNAL	43 :  STD_LOGIC;
SIGNAL	430 :  STD_LOGIC;
SIGNAL	431 :  STD_LOGIC;
SIGNAL	432 :  STD_LOGIC;
SIGNAL	433 :  STD_LOGIC;
SIGNAL	434 :  STD_LOGIC;
SIGNAL	435 :  STD_LOGIC;
SIGNAL	44 :  STD_LOGIC;
SIGNAL	440 :  STD_LOGIC;
SIGNAL	441 :  STD_LOGIC;
SIGNAL	442 :  STD_LOGIC;
SIGNAL	443 :  STD_LOGIC;
SIGNAL	444 :  STD_LOGIC;
SIGNAL	445 :  STD_LOGIC;
SIGNAL	45 :  STD_LOGIC;
SIGNAL	450 :  STD_LOGIC;
SIGNAL	451 :  STD_LOGIC;
SIGNAL	452 :  STD_LOGIC;
SIGNAL	453 :  STD_LOGIC;
SIGNAL	454 :  STD_LOGIC;
SIGNAL	455 :  STD_LOGIC;
SIGNAL	46 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	47 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	48 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	49 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	50 :  STD_LOGIC;
SIGNAL	500 :  STD_LOGIC;
SIGNAL	501 :  STD_LOGIC;
SIGNAL	502 :  STD_LOGIC;
SIGNAL	503 :  STD_LOGIC;
SIGNAL	504 :  STD_LOGIC;
SIGNAL	505 :  STD_LOGIC;
SIGNAL	51 :  STD_LOGIC;
SIGNAL	510 :  STD_LOGIC;
SIGNAL	511 :  STD_LOGIC;
SIGNAL	512 :  STD_LOGIC;
SIGNAL	513 :  STD_LOGIC;
SIGNAL	514 :  STD_LOGIC;
SIGNAL	515 :  STD_LOGIC;
SIGNAL	52 :  STD_LOGIC;
SIGNAL	53 :  STD_LOGIC;
SIGNAL	54 :  STD_LOGIC;
SIGNAL	55 :  STD_LOGIC;
SIGNAL	6 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	7 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	8 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	9 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	EMPTY_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	FF0_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF10_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF1_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF2_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF3_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF4_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF5_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF6_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF7_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF8_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FF9_OUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	FULL_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	HIGH :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	INIT :  STD_LOGIC;
SIGNAL	P_EN :  STD_LOGIC_VECTOR(51 DOWNTO 0);
SIGNAL	POP_ENABLE_INPUT :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	ZERO :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;

SIGNAL	GDFX_TEMP_SIGNAL_0 :  ARRAY2D0;

BEGIN 

GDFX_TEMP_SIGNAL_0 <= (515 & 514 & 513 & 512 & 511 & 510 & 505 & 504 & 503 & 502 & 501 & 500 & 49(5 DOWNTO 0) & 48(5 DOWNTO 0) & 47(5 DOWNTO 0) & 46(5 DOWNTO 0) & 455 & 454 & 453 & 452 & 451 & 450 & 445 & 444 & 443 & 442 & 441 & 440 & 435 & 434 & 433 & 432 & 431 & 430 & 425 & 424 & 423 & 422 & 421 & 420 & 415 & 414 & 413 & 412 & 411 & 410 & 405 & 404 & 403 & 402 & 401 & 400 & 39(5 DOWNTO 0) & 38(5 DOWNTO 0) & 37(5 DOWNTO 0) & 36(5 DOWNTO 0) & 355 & 354 & 353 & 352 & 351 & 350 & 345 & 344 & 343 & 342 & 341 & 340 & 335 & 334 & 333 & 332 & 331 & 330 & 325 & 324 & 323 & 322 & 321 & 320 & 315 & 314 & 313 & 312 & 311 & 310 & 305 & 304 & 303 & 302 & 301 & 300 & 29(5 DOWNTO 0) & 28(5 DOWNTO 0) & 27(5 DOWNTO 0) & 26(5 DOWNTO 0) & 255 & 254 & 253 & 252 & 251 & 250 & 245 & 244 & 243 & 242 & 241 & 240 & 235 & 234 & 233 & 232 & 231 & 230 & 225 & 224 & 223 & 222 & 221 & 220 & 215 & 214 & 213 & 212 & 211 & 210 & 205 & 204 & 203 & 202 & 201 & 200 & 19(5 DOWNTO 0) & 18(5 DOWNTO 0) & 17(5 DOWNTO 0) & 16(5 DOWNTO 0) & 155 & 154 & 153 & 152 & 151 & 150 & 145 & 144 & 143 & 142 & 141 & 140 & 135 & 134 & 133 & 132 & 131 & 130 & 125 & 124 & 123 & 122 & 121 & 120 & 115 & 114 & 113 & 112 & 111 & 110 & 105 & 104 & 103 & 102 & 101 & 100 & 9(5 DOWNTO 0) & 8(5 DOWNTO 0) & 7(5 DOWNTO 0) & 6(5 DOWNTO 0) & 55 & 54 & 53 & 52 & 51 & 50 & 45 & 44 & 43 & 42 & 41 & 40 & 35 & 34 & 33 & 32 & 31 & 30 & 25 & 24 & 23 & 22 & 21 & 20 & 15 & 14 & 13 & 12 & 11 & 10 & 0(5 DOWNTO 0));


b2v_counter : lpm_counter0
PORT MAP(sclr => RST,
		 sload => EMPTY_ALTERA_SYNTHESIZED,
		 sset => INIT,
		 updown => SYNTHESIZED_WIRE_0,
		 clock => CLK,
		 cnt_en => SYNTHESIZED_WIRE_1,
		 data => ZERO,
		 q => NUM);


b2v_inst : lpm_ff_0
PORT MAP(enable => P_EN(0),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_2,
		 q => FF0_OUT);


b2v_inst1 : lpm_mux2
PORT MAP(data0x => ADDR,
		 data1x => ZERO,
		 data2x => HIGH,
		 data3x => HIGH,
		 sel => MODE,
		 result => POP_ENABLE_INPUT);


POP <= ENABLE AND MODE(1) AND MODE(0) AND SYNTHESIZED_WIRE_3;


b2v_inst11 : lpm_ff_1
PORT MAP(enable => P_EN(1),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_4,
		 q => FF1_OUT);


SYNTHESIZED_WIRE_3 <= NOT(FULL_ALTERA_SYNTHESIZED);



b2v_inst13 : g27_pop_enable
PORT MAP(clk => CLK,
		 N => POP_ENABLE_INPUT,
		 P_EN => P_EN);


INIT <= SYNTHESIZED_WIRE_5 AND MODE(0);


SYNTHESIZED_WIRE_5 <= NOT(MODE(1));



b2v_inst16 : lpm_ff_2
PORT MAP(enable => P_EN(7),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_6,
		 q => FF7_OUT);



b2v_inst18 : lpm_ff_3
PORT MAP(enable => P_EN(2),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_7,
		 q => FF2_OUT);



b2v_inst2 : busmux_4
PORT MAP(sel => MODE(0),
		 dataa => DATA,
		 datab => FF1_OUT,
		 result => SYNTHESIZED_WIRE_2);


b2v_inst20 : lpm_ff_5
PORT MAP(enable => P_EN(4),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_8,
		 q => FF4_OUT);



b2v_inst22 : lpm_mux_6
PORT MAP(data => GDFX_TEMP_SIGNAL_0,
		 sel => ADDR);


b2v_inst23 : lpm_ff_7
PORT MAP(enable => P_EN(6),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_9,
		 q => FF6_OUT);


b2v_inst24 : busmux_8
PORT MAP(sel => MODE(0),
		 dataa => FF4_OUT,
		 datab => FF6_OUT,
		 result => SYNTHESIZED_WIRE_11);


b2v_inst25 : busmux_9
PORT MAP(sel => MODE(0),
		 dataa => FF6_OUT,
		 datab => FF8_OUT,
		 result => SYNTHESIZED_WIRE_6);


SYNTHESIZED_WIRE_0 <= NOT(MODE(0));



SYNTHESIZED_WIRE_1 <= MODE(1) AND SYNTHESIZED_WIRE_10;


b2v_inst28 : busmux_10
PORT MAP(sel => MODE(0),
		 dataa => FF5_OUT,
		 datab => FF7_OUT,
		 result => SYNTHESIZED_WIRE_9);


SYNTHESIZED_WIRE_10 <= NOT(FULL_ALTERA_SYNTHESIZED);



b2v_inst3 : busmux_11
PORT MAP(sel => MODE(0),
		 dataa => FF0_OUT,
		 datab => FF2_OUT,
		 result => SYNTHESIZED_WIRE_4);


b2v_inst30 : lpm_ff_12
PORT MAP(enable => P_EN(5),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_11,
		 q => FF5_OUT);


b2v_inst31 : busmux_13
PORT MAP(sel => MODE(0),
		 dataa => FF7_OUT,
		 datab => FF9_OUT,
		 result => SYNTHESIZED_WIRE_12);


b2v_inst32 : lpm_ff_14
PORT MAP(enable => P_EN(8),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_12,
		 q => FF8_OUT);


b2v_inst33 : busmux_15
PORT MAP(sel => MODE(0),
		 dataa => FF8_OUT,
		 datab => FF10_OUT,
		 result => SYNTHESIZED_WIRE_13);


b2v_inst34 : lpm_ff_16
PORT MAP(enable => P_EN(9),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_13,
		 q => FF9_OUT);


b2v_inst35 : busmux_17
PORT MAP(sel => MODE(0),
		 dataa => FF9_OUT,
		 datab => ZERO,
		 result => SYNTHESIZED_WIRE_14);


b2v_inst37 : lpm_ff_18
PORT MAP(enable => P_EN(10),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_14,
		 q => FF10_OUT);


b2v_inst4 : busmux_19
PORT MAP(sel => MODE(0),
		 dataa => FF2_OUT,
		 datab => FF4_OUT,
		 result => SYNTHESIZED_WIRE_15);


b2v_inst5 : lpm_ff_20
PORT MAP(enable => P_EN(3),
		 clock => CLK,
		 sset => INIT,
		 sclr => RST,
		 data => SYNTHESIZED_WIRE_15,
		 q => FF3_OUT);


b2v_inst6 : busmux_21
PORT MAP(sel => MODE(0),
		 dataa => FF1_OUT,
		 datab => FF3_OUT,
		 result => SYNTHESIZED_WIRE_7);


SYNTHESIZED_WIRE_16 <= NOT(MODE(0));



PUSH <= ENABLE AND MODE(1) AND SYNTHESIZED_WIRE_16 AND SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_17 <= NOT(FULL_ALTERA_SYNTHESIZED);



b2v_mux4 : busmux_22
PORT MAP(sel => MODE(0),
		 dataa => FF3_OUT,
		 datab => FF5_OUT,
		 result => SYNTHESIZED_WIRE_8);

EMPTY <= EMPTY_ALTERA_SYNTHESIZED;
FULL <= FULL_ALTERA_SYNTHESIZED;

FULL_ALTERA_SYNTHESIZED <= '0';
HIGH <= "111111";
ZERO <= "000000";
END bdf_type;