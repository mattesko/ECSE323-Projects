library verilog;
use verilog.vl_types.all;
entity g27_8bit_adder_vlg_vec_tst is
end g27_8bit_adder_vlg_vec_tst;
