library verilog;
use verilog.vl_types.all;
entity deal_schematic_vlg_vec_tst is
end deal_schematic_vlg_vec_tst;
