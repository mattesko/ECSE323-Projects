library verilog;
use verilog.vl_types.all;
entity testing_vlg_vec_tst is
end testing_vlg_vec_tst;
