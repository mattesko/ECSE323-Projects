library verilog;
use verilog.vl_types.all;
entity g27_Modulo_13 is
    port(
        O               : out    vl_logic_vector(3 downto 0);
        \IN\            : in     vl_logic_vector(5 downto 0)
    );
end g27_Modulo_13;
